library ieee;
use ieee.std_logic_1164.all;

library work;
use work.proj.all;

entity test_project__tpch__const_date_generator_s_com is
  port (
    clk : in std_logic;
    rst : in std_logic;
    date_output_valid : out std_logic;
    date_output_ready : in std_logic;
    date_output_data : out std_logic_vector(25 downto 0);
    date_output_last : out std_logic;
    date_output_strb : out std_logic
  );
end test_project__tpch__const_date_generator_s_com;

architecture Behavioral of test_project__tpch__const_date_generator_s_com is
begin
end Behavioral;